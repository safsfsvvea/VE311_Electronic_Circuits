** Profile: "SCHEMATIC1-sim3_2"  [ D:\pspice\hw3\hw3_2-pspicefiles\schematic1\sim3_2.sim ] 

** Creating circuit file "sim3_2.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../hw3_2-pspicefiles/hw3_2.lib" 
* From [PSPICE NETLIST] section of C:\Users\ZWK\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.DC LIN V_V3 0.45V 0.55V 0.0001 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
